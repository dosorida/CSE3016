`timescale 1ns / 1ps

module binary_counter_tb;

reg clk, rst;
wire[1:0] out;

binary_counter u_binary_counter (
.clk (clk ),
.rst (rst ),
.out (out )
);

always #10 clk = ~clk;

initial begin
clk = 1'b0;
rst = 1'b0;
#20 rst <= 1'b1;
#80 rst <= 1'b0;
#50 rst <= 1'b1;
end  

initial begin 
    #1000
    $finish;
end

endmodule
