`timescale 1ns / 1ps
module buff(
input a,
output y
);
assign y=a;
endmodule